    `timescale 1ns / 1ps
    
    module SPMemory(input clk,input sclk,input[31:0] addr,input MemRead, input MemWrite,
     input [2:0]func3,input [31:0]readData2,output reg  [31:0]  data_out);
      reg [7:0] mem [(1024-1):0]; 
    
    //***************instruction memory***********//
    always @(*)
    begin
    if (sclk)
     data_out ={ mem[addr+3],mem[addr+2],mem[addr+1],mem[addr+0]};
     else  if ( func3 == 3'b010)//\\lw
          data_out = MemRead ? { mem[1024/2+addr+3],mem[1024/2+addr+2]
          ,mem[1024/2+addr+1],mem[1024/2+addr+0]}:0;
     else if( func3 == 3'b000)//lb
           data_out = MemRead ? mem[1024/2+addr+0]:0;
     else if ( func3 == 3'b001)//Lh
           data_out = MemRead ? { 
           mem[1024/2+addr+1],mem[1024/2+addr+0]}:0;
     else if ( func3 == 3'b100)
           data_out = MemRead ? {24'h0,mem[1024/2+addr+0]}:0;
     else if ( func3 == 3'b101)
            data_out = MemRead ? { 16'h0,
            mem[1024/2+addr+1],mem[1024/2+addr+0]}:0;
    
       end
    
    initial begin
    
    // R_type
    //{mem[3],mem[2],mem[1],mem[0]}=32'b00000000000000000000000000110011;//NOP 
    //{mem[7],mem[6],mem[5],mem[4]}=32'b00000000000000000010001010000011;
    //{mem[11],mem[10],mem[9],mem[8]}=32'b00000000010000000010001100000011;
    //{mem[15],mem[14],mem[13],mem[12]}=32'b00000000100000000010001110000011;
    //{mem[19],mem[18],mem[17],mem[16]}=32'b00000000010100110000111000110011;
    //{mem[23],mem[22],mem[21],mem[20]}=32'b01000000010100110000111010110011;
    //{mem[27],mem[26],mem[25],mem[24]}=32'b00000000010100110111111100110011;
    //{mem[31],mem[30],mem[29],mem[28]}=32'b00000000010100110100111110110011;
    
    // I_TYPE completed test
    //{mem[7],mem[6],mem[5],mem[4]}=32'b00000000010000000010001100000011; 
    //{mem[11],mem[10],mem[9],mem[8]}=32'b00000000101000110000111000010011;
    //{mem[15],mem[14],mem[13],mem[12]}=32'b00000000101000110111111100010011;
    //{mem[19],mem[18],mem[17],mem[16]}=32'b00000000101000110100111110010011;
    //{mem[23],mem[22],mem[21],mem[20]}=32'b00000000101000110110010000010011;
    //{mem[27],mem[26],mem[25],mem[24]}=32'b00000000001000110001010010010011;
    //{mem[31],mem[30],mem[29],mem[28]}=32'b00000000101000110010100100010011;
    //{mem[35],mem[34],mem[33],mem[32]}=32'b00000000101000110011100110010011;
    //{mem[39],mem[38],mem[37],mem[36]}=32'b01000000001000110101101000010011;
    //{mem[43],mem[42],mem[41],mem[40]}=32'b00000000101000110101101010010011;
    
    //Jal_Auipc_lui
    //{mem[7],mem[6],mem[5],mem[4]}=32'b00000000000000000010001100000011;
    //{mem[11],mem[10],mem[9],mem[8]}=32'b00000000010000000010001110000011;
    //{mem[15],mem[14],mem[13],mem[12]}=32'b00000000100000000010111000000011;
    //{mem[19],mem[18],mem[17],mem[16]}=32'b00000000100000000000000011101111;
    //{mem[23],mem[22],mem[21],mem[20]}=32'b00000000000100110000001100010011;
    //{mem[27],mem[26],mem[25],mem[24]}=32'b00000010011100010000001110010111;
    //{mem[31],mem[30],mem[29],mem[28]}=32'b00000010011100010000111000110111;
    //{mem[35],mem[34],mem[33],mem[32]}=32'b00000000000000000000111010010011;
    //{mem[39],mem[38],mem[37],mem[36]}=32'b00000010010011101000001011100111;
    //{mem[43],mem[42],mem[41],mem[40]}=32'b00000000000100110000001100010011;
    //{mem[46],mem[45],mem[44],mem[44]}=32'b00000001110000000010011000100011;
    
    
    //lab progeam to test the hards
    //{mem[7],mem[6],mem[5],mem[4]}=32'b000000000000_00000_010_00001_0000011 ;
    // {mem[11],mem[10],mem[9],mem[8]}=32'b000000000100_00000_010_00010_0000011 ; 
    //{mem[15],mem[14],mem[13],mem[12]}=32'b000000001000_00000_010_00011_0000011 ; 
    //{mem[19],mem[18],mem[17],mem[16]}=32'b0000000_00010_00001_110_00100_0110011 ;
    //{mem[23],mem[22],mem[21],mem[20]}=32'b0_000000_00011_00100_000_0100_0_1100011 ;
    // {mem[27],mem[26],mem[25],mem[24]}=32'b0000000_00010_00001_000_00011_0110011 ; 
    //{mem[31],mem[30],mem[29],mem[28]}=32'b0000000_00010_00011_000_00101_0110011 ; 
    //{mem[35],mem[34],mem[33],mem[32]}=32'b0000000_00101_00000_010_01100_0100011; 
    //{mem[39],mem[38],mem[37],mem[36]}=32'b000000001100_00000_010_00110_0000011 ; 
    //{mem[43],mem[42],mem[41],mem[40]}=32'b0000000_00001_00110_111_00111_0110011 ;
    //{mem[47],mem[46],mem[45],mem[44]}=32'b0100000_00010_00001_000_01000_0110011 ;
    //{mem[51],mem[50],mem[49],mem[48]}=32'b0000000_00010_00001_000_00000_0110011 ;
    //{mem[55],mem[54],mem[53],mem[52]}=32'b0000000_00001_00000_000_01001_0110011;
    
    
       
        $readmemh("./test_all_instructions.mem", mem);

//$readmemh("./jalr_jal.mem", mem);
    
    end
    
    
    
    
    
    
    
    //mem[6]=32'b00000000010100110100111110110011;
    //mem[7]=32'b00000000010100110110010000110011;
    //mem[8]=32'b00000000011100110001010010110011;
    //mem[9]=32'b00000000010100110010100100110011;
    //mem[10]=32'b00000000010100110011100110110011;
    //mem[11]=32'b01000000011100110101101000110011;
    //mem[12]=32'b00000000010100110101101010110011
    
    
    //mem[7]=32'b00000001110000000010011000100011;
    //mem[8]=32'b00000000000000000000000001110011;
    //**********data memory*************//
    always @(posedge clk)
    begin
    if (MemWrite==1 && func3 ==3'b010)
    { mem[1024/2+addr+3],mem[1024/2+addr+2]
    ,mem[1024/2+addr+1],mem[1024/2+addr+0]} <= readData2[31:0];
      
      else if (MemWrite==1 && func3 ==3'b000)//sb
      mem[1024/2+addr+0] <= {readData2[7:0]};
      else if (MemWrite==1 && func3 ==3'b001)//sh
      {  mem[1024/2+addr+1],mem[1024/2+addr+0]} <= readData2[15:0];
      
      
      end
      
    //  always @(*)
    //  begin
      
    //   if ( func3 == 3'b010)//\\lw
    //      data_out = MemRead ? { mem[2*1024+addr+3],mem[2*1024+addr+2]
    //      ,mem[2*1024+addr+1],mem[2*1024+addr+0]}:0;
    //        else if( func3 == 3'b000)//lb
    //         data_out = MemRead ? mem[2*1024+addr+0]:0;
    //         else if ( func3 == 3'b001)//Lh
    //          data_out = MemRead ? { 
    //          mem[2*1024+addr+1],mem[2*1024+addr+0]}:0;
    //           else if ( func3 == 3'b100)
    //           data_out = MemRead ? {24'h0,mem[2*1024+addr+0]}:0;
    //            else if ( func3 == 3'b101)
    //              data_out = MemRead ? { 16'h0,
    //            mem[2*1024+addr+1],mem[2*1024+addr+0]}:0;
               
    //    end
        //store
        
      
       
    
    
    
    initial
     begin
     {mem[1024/2+3],mem[1024/2+2],mem[1024/2+1],mem[1024/2+0]}=32'd17;
     {mem[1024/2+7],mem[1024/2+6],mem[1024/2+5],mem[1024/2+4]}=32'd9;
     {mem[1024/2+11],mem[1024/2+10],mem[1024/2+9],mem[1024/2+8]}=32'd25;
      {mem[1024/2+19],mem[1024/2+18],mem[1024/2+17],mem[1024/2+16]}=32'd100000000;
     end
    
    
    
     
     
     
    
    
    
    
    
    
    
    
    
    
    
    
    endmodule
